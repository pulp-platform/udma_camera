package cpi_pkg;
	 // cpi structure
	typedef struct packed{
		logic pclk_i;
		logic hsync_i;
		logic vsync_i;
		logic data0_i;
		logic data1_i;
		logic data2_i;
		logic data3_i;
		logic data4_i;
		logic data5_i;
		logic data6_i;
		logic data7_i;
	}pad_to_cpi_t;
endpackage