package camera_verisuite_pkg;
	typedef struct packed {
		logic [31:0] value;
		logic [31:0] addr;
	}cfg_reg_t;
endpackage